library verilog;
use verilog.vl_types.all;
entity example_verilog_vlg_vec_tst is
end example_verilog_vlg_vec_tst;
